module tb_Register();




endmodule 